module mem(input  logic        clk, we,
           input  logic [31:0] a, wd,
           output logic [31:0] rd);

  logic  [31:0] RAM[63:0]; // 64 addresses of one word (32 bits)

  // initialize memory with instructions
  initial
    begin
      $readmemh("memfile.dat",RAM);  // Instructions are in hexadecimal.  Load the program.
                                     
    end

  assign rd = RAM[a[31:2]]; // word

  always_ff @(posedge clk)
    if (we)
      RAM[a[31:2]] <= wd; // Only write on enable
endmodule